----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    12:07:50 05/11/2018 
-- Design Name: 
-- Module Name:    pixelBuffer - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity pixelBuffer is
    Port ( iWR_CLK : in  STD_LOGIC;
			  iRD_CLK : in STD_LOGIC;
           inRST : in  STD_LOGIC;
           oCMD_EN : out  STD_LOGIC;
           oCMD_INSTR : out  STD_LOGIC_VECTOR (2 downto 0);
           oCMD_BL : out  STD_LOGIC_VECTOR (5 downto 0);
           oCMD_BYTE_ADDR : out  STD_LOGIC_VECTOR (29 downto 0);
           iCMD_EMPTY : in  STD_LOGIC;
           iCMD_FULL : in  STD_LOGIC;
           oRD_EN : out  STD_LOGIC;
           iRD_DATA : in  STD_LOGIC_VECTOR (31 downto 0);
           iRD_FULL : in  STD_LOGIC;
           iRD_EMPTY : in  STD_LOGIC;
           iRD_OVERFLOW : in  STD_LOGIC;
           iRD_ERROR : in  STD_LOGIC;
           iRD_COUNT : in  STD_LOGIC_VECTOR (6 downto 0);
			  iFIFO_RD_EN : in STD_LOGIC;
			  iSTART : in STD_LOGIC;
			  oRGB : out STD_LOGIC_VECTOR (23 downto 0));
end pixelBuffer;

architecture Behavioral of pixelBuffer is

	type tREAD_STATE is (IDLE, SET_CMD, WAIT_DATA, READ_DATA, CHECK_FIFO, WAIT_FIFO);
	signal sSTATE, sNEXT_STATE : tREAD_STATE;

	signal sINV_RST : STD_LOGIC;
	signal sFIFO_FULL : STD_LOGIC;
	signal sFIFO_EMPTY : STD_LOGIC;
	signal sFIFO_RD_EN : STD_LOGIC;
	signal sFIFO_WR_EN : STD_LOGIC;
	signal sPOS_X : STD_LOGIC_VECTOR(10 downto 0);
	signal sPOS_Y : STD_LOGIC_VECTOR(9 downto 0);
	signal sPOS_WE : STD_LOGIC;
	signal sCOMBINED_EN : STD_LOGIC;
	
begin
	
	sINV_RST <= not inRST;	
		
	oCMD_INSTR <= "001";
	oCMD_BL <= (others => '1');
	oCMD_BYTE_ADDR <= "000000" & sPOS_Y & "00" & sPOS_X(9 downto 0) & "00";
		
	sCOMBINED_EN <= sFIFO_RD_EN and iFIFO_RD_EN;
		
	process(iRD_CLK, inRST) begin
		if(inRST = '0') then
			sFIFO_RD_EN <= '0';
		elsif(iRD_CLK'event and iRD_CLK = '1') then
			if(sFIFO_FULL = '1' and iSTART = '1' and sFIFO_EMPTY = '0') then
				sFIFO_RD_EN <= '1';
			end if;
		end if;
	end process;
	
	process(iWR_CLK, inRST) begin
		if(inRST = '0') then
			sPOS_X <= (others => '0');
			sPOS_Y <= (others => '0');
		elsif(iWR_CLK'event and iWR_CLK = '1') then
			if(sPOS_WE = '1') then
				if(sPOS_X = 960) then
					sPOS_X <= (others => '0');
					if(sPOS_Y = 767) then
						sPOS_Y <= (others => '0');
					else
						sPOS_Y <= sPOS_Y + 1;
					end if;
				else
					sPOS_X <= sPOS_X + 64;
				end if;
			end if;
		end if;
	end process;
		
	process(iWR_CLK, inRST) begin
		if(inRST = '0') then
			sSTATE <= IDLE;
		elsif(iWR_CLK'event and iWR_CLK = '1') then
			sSTATE <= sNEXT_STATE;
		end if;
	end process;
	
	process(sSTATE, iRD_FULL, iRD_COUNT, sFIFO_FULL) begin
		case sSTATE is
			when IDLE =>
					sNEXT_STATE <= SET_CMD;
			when SET_CMD =>
				sNEXT_STATE <= WAIT_DATA;
			when WAIT_DATA =>
				if(iRD_FULL = '1') then
					sNEXT_STATE <= READ_DATA;
				else
					sNEXT_STATE <= WAIT_DATA;
				end if;
			when READ_DATA =>
				if(iRD_COUNT = 1) then
					sNEXT_STATE <= CHECK_FIFO;
				else
					sNEXT_STATE <= READ_DATA;
				end if;
			when CHECK_FIFO =>
				if(sFIFO_FULL = '1') then
					sNEXT_STATE <= WAIT_FIFO;
				else
					sNEXT_STATE <= SET_CMD;
				end if;
			when others =>
				if(sFIFO_FULL = '0') then
					sNEXT_STATE <= SET_CMD;
				else
					sNEXT_STATE <= WAIT_FIFO;
				end if;
		end case;
	end process;
	
	process(sSTATE) begin
		case sSTATE is
			when IDLE =>
				oCMD_EN <= '0';
				oRD_EN <= '0';
				sPOS_WE <= '0';
				sFIFO_WR_EN <= '0';
				
			when SET_CMD =>
				oCMD_EN <= '1';
				oRD_EN <= '0';
				sPOS_WE <= '1';
				sFIFO_WR_EN <= '0';
			
			when WAIT_DATA =>
				oCMD_EN <= '0';
				oRD_EN <= '0';
				sPOS_WE <= '0';
				sFIFO_WR_EN <= '0';
				
			when READ_DATA =>
				oCMD_EN <= '0';
				oRD_EN <= '1';
				sPOS_WE <= '0';
				sFIFO_WR_EN <= '1';
				
			when others =>
				oCMD_EN <= '0';
				oRD_EN <= '0';
				sPOS_WE <= '0';
				sFIFO_WR_EN <= '0';
				
		end case;
	end process;
	
	fifo : entity work.fif0
		port map(
		 rst => sINV_RST,
		 wr_clk => iWR_CLK,
		 rd_clk => iRD_CLK,
		 din => iRD_DATA(23 downto 0),
		 wr_en => sFIFO_WR_EN,
		 rd_en => sCOMBINED_EN,
		 dout => oRGB,
		 full => open,
		 empty => sFIFO_EMPTY,
		 prog_full => sFIFO_FULL
  );
  
  
end Behavioral;

